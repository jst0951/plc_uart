library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_arith.all;
  use ieee.std_logic_unsigned.all;
  
entity tb_plc_uart is end;

architecture BEH of tb_plc_uart is
  
  component plc_uart is
  port(
    nRst  : in std_logic;
    clk   : in std_logic;
    -- PLC INPUT
    Y20   : in std_logic;
    Y21   : in std_logic;
    -- UART TX BUSY
    busy  : in std_logic;
    -- UART TX OUTPUT
    tx_data  : out std_logic_vector(7 downto 0);
    start_sig : out std_logic
  );
  end component;
  
  component uart_tx is
  port(
    nRst  : in std_logic;
    clk   : in std_logic;
    start_sig : in std_logic;
    data      : in std_logic_vector(7 downto 0);
    tx        : out std_logic;
    busy      : out std_logic
  );
  end component;
  
  -- common
  signal nRst : std_logic;
  signal clk  : std_logic;
  -- plc_uart
  signal Y20 : std_logic;
  signal Y21 : std_logic;
  -- uart_tx
  signal tx_data : std_logic_vector(7 downto 0);
  signal start_sig : std_logic;
  signal tx : std_logic;
  signal busy : std_logic;
  -- internal counter
  signal int_cnt : std_logic_vector(99 downto 0);
  
begin
  U_plc_uart : plc_uart
  port map(
    nRst  => nRst,
    clk   => clk,
    Y20   => Y20,
    Y21   => Y21,
    busy  => busy,
    tx_data => tx_data,
    start_sig => start_sig
  );
  
  U_uart_tx : uart_tx
  port map(
    nRst  => nRst,
    clk   => clk,
    start_sig => start_sig,
    data      => tx_data,
    tx    => tx,
    busy  => busy
  );
  
  -- nRst
  process
  begin
    nRst <= '0', '1' after 200 ns;
    wait for 1 sec;
  end process;
  
  -- clk
  process
  begin
    clk <= '0', '1' after 5 ns;
    wait for 10 ns;
  end process;
  
  -- cylinder input setting
  process(nRSt, clk)
  begin
    if(nRst = '0') then
      int_cnt <= (others => '0');
    elsif rising_edge(clk) then
      int_cnt <= int_cnt + 1;
    end if;
  end process;
  Y20 <= '1' when 100 < int_cnt and int_cnt < 200 else '0';
  Y21 <= '1' when 200100 < int_cnt and int_cnt < 200200 else '0';
end BEH;